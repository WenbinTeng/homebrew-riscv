module _74x154 (
    input [3:0] a,  // Address Inputs
    input [1:0] g,  // Enable (Active LOW) Inputs
    output [15:0] o // Active LOW Outputs
);

    reg [15:0] out;

    always @(*) begin
        case (a)
            4'b0000: out = 16'b1111111111111110;
            4'b0001: out = 16'b1111111111111101;
            4'b0010: out = 16'b1111111111111011;
            4'b0011: out = 16'b1111111111110111;
            4'b0100: out = 16'b1111111111101111;
            4'b0101: out = 16'b1111111111011111;
            4'b0110: out = 16'b1111111110111111;
            4'b0111: out = 16'b1111111101111111;
            4'b1000: out = 16'b1111111011111111;
            4'b1001: out = 16'b1111110111111111;
            4'b1010: out = 16'b1111101111111111;
            4'b1011: out = 16'b1111011111111111;
            4'b1100: out = 16'b1110111111111111;
            4'b1101: out = 16'b1101111111111111;
            4'b1110: out = 16'b1011111111111111;
            4'b1111: out = 16'b0111111111111111;
        endcase
    end

    assign o = !g[1] & !g[0] ? out : 16'b1111111111111111;
    
endmodule